import FIFO::*;
import FIFOF::*;
import Clocks::*;
import Vector::*;

import BRAM::*;
import BRAMFIFO::*;

import PageSorter::*;

interface DRAMMergerIfc;
endinterface


module mkDRAMMerger (DRAMMergerIfc);
endmodule
