module null_reset_n ( RESET_N );
	output RESET_N;
	assign RESET_N = 1;
endmodule
